# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__a211oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.350000 3.855000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.300000 6.115000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.894000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 7.555000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.685800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.570000 0.785000 3.760000 0.960000 ;
        RECT 2.570000 0.960000 6.490000 1.010000 ;
        RECT 2.570000 1.010000 8.515000 1.130000 ;
        RECT 5.380000 0.350000 5.630000 0.960000 ;
        RECT 6.320000 0.350000 6.490000 0.960000 ;
        RECT 6.320000 1.130000 8.515000 1.180000 ;
        RECT 6.795000 1.950000 7.895000 2.120000 ;
        RECT 6.795000 2.120000 6.965000 2.735000 ;
        RECT 7.180000 0.350000 8.515000 1.010000 ;
        RECT 7.695000 2.120000 7.895000 2.735000 ;
        RECT 7.725000 1.180000 8.515000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.345000  1.950000 6.145000 2.120000 ;
      RECT 0.345000  2.120000 0.675000 2.980000 ;
      RECT 0.420000  0.350000 0.670000 1.010000 ;
      RECT 0.420000  1.010000 2.390000 1.180000 ;
      RECT 0.850000  0.085000 1.180000 0.840000 ;
      RECT 0.875000  2.290000 1.045000 3.245000 ;
      RECT 1.245000  2.120000 1.495000 2.980000 ;
      RECT 1.360000  0.350000 1.530000 1.010000 ;
      RECT 1.695000  2.290000 2.025000 3.245000 ;
      RECT 1.710000  0.085000 2.040000 0.840000 ;
      RECT 2.220000  0.350000 4.190000 0.615000 ;
      RECT 2.220000  0.615000 2.390000 1.010000 ;
      RECT 2.225000  2.120000 2.395000 2.980000 ;
      RECT 2.595000  2.290000 2.925000 3.245000 ;
      RECT 3.125000  2.120000 3.295000 2.980000 ;
      RECT 3.495000  2.290000 3.825000 3.245000 ;
      RECT 4.025000  1.820000 4.275000 1.950000 ;
      RECT 4.025000  2.120000 4.275000 2.980000 ;
      RECT 4.465000  2.290000 4.795000 2.905000 ;
      RECT 4.465000  2.905000 8.395000 3.075000 ;
      RECT 4.995000  2.120000 5.165000 2.735000 ;
      RECT 5.365000  2.290000 5.695000 2.905000 ;
      RECT 5.810000  0.085000 6.140000 0.790000 ;
      RECT 5.895000  2.120000 6.145000 2.735000 ;
      RECT 6.315000  1.950000 6.595000 2.905000 ;
      RECT 6.670000  0.085000 7.000000 0.840000 ;
      RECT 7.165000  2.290000 7.495000 2.905000 ;
      RECT 8.065000  2.120000 8.395000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ls__a211oi_4
END LIBRARY
