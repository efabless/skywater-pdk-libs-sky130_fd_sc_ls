# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__nor4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 1.180000 3.715000 1.540000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.285000 1.320000 2.625000 1.650000 ;
        RECT 2.455000 1.650000 2.625000 1.710000 ;
        RECT 2.455000 1.710000 4.215000 1.880000 ;
        RECT 3.885000 0.280000 4.215000 1.710000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.170000 0.700000 1.320000 ;
        RECT 0.425000 1.320000 2.075000 1.500000 ;
        RECT 1.565000 1.500000 2.075000 1.650000 ;
        RECT 1.565000 1.650000 1.795000 2.150000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.447000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.330000 0.435000 0.660000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.808000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.830000 1.880000 0.980000 ;
        RECT 0.085000 0.980000 2.880000 1.000000 ;
        RECT 0.085000 1.000000 0.255000 1.670000 ;
        RECT 0.085000 1.670000 1.385000 1.840000 ;
        RECT 0.615000 1.840000 1.385000 2.150000 ;
        RECT 1.550000 0.350000 1.880000 0.830000 ;
        RECT 1.550000 1.000000 2.880000 1.150000 ;
        RECT 2.550000 0.350000 2.880000 0.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  2.010000 0.445000 2.320000 ;
      RECT 0.115000  2.320000 2.285000 2.490000 ;
      RECT 0.115000  2.490000 0.365000 3.000000 ;
      RECT 0.565000  2.660000 1.835000 2.980000 ;
      RECT 0.605000  0.085000 1.380000 0.600000 ;
      RECT 2.035000  1.820000 2.285000 2.050000 ;
      RECT 2.035000  2.050000 4.205000 2.220000 ;
      RECT 2.035000  2.220000 2.285000 2.320000 ;
      RECT 2.035000  2.490000 2.285000 2.980000 ;
      RECT 2.050000  0.085000 2.380000 0.810000 ;
      RECT 2.475000  2.390000 3.755000 2.560000 ;
      RECT 2.475000  2.560000 2.805000 3.000000 ;
      RECT 2.975000  2.730000 3.305000 3.245000 ;
      RECT 3.050000  0.085000 3.380000 1.010000 ;
      RECT 3.505000  2.560000 3.755000 3.000000 ;
      RECT 3.940000  2.220000 4.205000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ls__nor4_2
END LIBRARY
