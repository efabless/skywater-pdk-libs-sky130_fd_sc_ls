# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__o22ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.910000 1.350000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665000 1.300000 3.335000 1.390000 ;
        RECT 2.665000 1.390000 3.715000 1.630000 ;
        RECT 3.485000 1.630000 3.715000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.350000 1.815000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.212200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 0.595000 0.945000 1.010000 ;
        RECT 0.615000 1.010000 2.275000 1.180000 ;
        RECT 1.570000 1.950000 3.310000 1.970000 ;
        RECT 1.570000 1.970000 2.275000 2.120000 ;
        RECT 1.570000 2.120000 1.800000 2.735000 ;
        RECT 1.615000 0.595000 1.945000 1.010000 ;
        RECT 2.045000 1.180000 2.275000 1.800000 ;
        RECT 2.045000 1.800000 3.310000 1.950000 ;
        RECT 3.060000 1.970000 3.310000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.255000 2.785000 0.425000 ;
      RECT 0.115000  0.425000 0.445000 1.130000 ;
      RECT 0.120000  1.950000 1.400000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.570000  2.290000 0.900000 3.245000 ;
      RECT 1.070000  2.120000 1.400000 2.905000 ;
      RECT 1.070000  2.905000 2.300000 3.075000 ;
      RECT 1.115000  0.425000 1.445000 0.840000 ;
      RECT 1.970000  2.290000 2.300000 2.905000 ;
      RECT 2.115000  0.425000 2.785000 0.840000 ;
      RECT 2.455000  0.840000 2.785000 0.960000 ;
      RECT 2.455000  0.960000 3.755000 1.010000 ;
      RECT 2.455000  1.010000 4.685000 1.130000 ;
      RECT 2.530000  2.140000 2.860000 2.905000 ;
      RECT 2.530000  2.905000 3.680000 3.075000 ;
      RECT 2.955000  0.085000 3.285000 0.790000 ;
      RECT 3.505000  0.350000 3.755000 0.960000 ;
      RECT 3.505000  1.130000 4.685000 1.180000 ;
      RECT 3.510000  1.950000 4.660000 2.120000 ;
      RECT 3.510000  2.120000 3.680000 2.905000 ;
      RECT 3.880000  2.290000 4.130000 3.245000 ;
      RECT 3.925000  0.085000 4.255000 0.840000 ;
      RECT 4.330000  2.120000 4.660000 2.980000 ;
      RECT 4.435000  0.350000 4.685000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ls__o22ai_2
END LIBRARY
