# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__dlrbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.260000 0.805000 1.930000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.260000 1.820000 6.590000 2.070000 ;
        RECT 6.285000 0.770000 6.615000 1.130000 ;
        RECT 6.285000 1.130000 6.455000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.572800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.205000 0.880000 8.575000 1.050000 ;
        RECT 8.225000 1.820000 8.575000 2.980000 ;
        RECT 8.405000 1.050000 8.575000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.570000 1.180000 6.115000 1.550000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.237000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.260000 1.285000 1.930000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.085000  0.540000 0.445000 1.090000 ;
      RECT 0.085000  1.090000 0.255000 2.100000 ;
      RECT 0.085000  2.100000 1.155000 2.270000 ;
      RECT 0.085000  2.270000 0.445000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 1.090000 ;
      RECT 0.645000  2.440000 0.815000 3.245000 ;
      RECT 0.985000  2.270000 1.155000 2.650000 ;
      RECT 0.985000  2.650000 1.965000 2.820000 ;
      RECT 1.125000  0.350000 1.625000 1.090000 ;
      RECT 1.325000  2.100000 1.625000 2.140000 ;
      RECT 1.325000  2.140000 2.475000 2.310000 ;
      RECT 1.325000  2.310000 1.625000 2.480000 ;
      RECT 1.455000  1.090000 1.625000 2.100000 ;
      RECT 1.795000  0.350000 2.125000 0.780000 ;
      RECT 1.795000  0.780000 3.885000 0.950000 ;
      RECT 1.795000  0.950000 2.125000 0.960000 ;
      RECT 1.795000  0.960000 1.965000 1.720000 ;
      RECT 1.795000  1.720000 2.135000 1.970000 ;
      RECT 1.795000  2.480000 2.830000 2.650000 ;
      RECT 2.135000  1.130000 3.530000 1.300000 ;
      RECT 2.135000  1.300000 2.475000 1.550000 ;
      RECT 2.295000  0.085000 2.835000 0.600000 ;
      RECT 2.305000  1.550000 2.475000 2.140000 ;
      RECT 2.425000  2.820000 2.755000 3.245000 ;
      RECT 2.660000  1.470000 2.985000 1.800000 ;
      RECT 2.660000  1.800000 2.830000 2.480000 ;
      RECT 3.010000  1.970000 3.325000 2.140000 ;
      RECT 3.010000  2.140000 3.180000 2.905000 ;
      RECT 3.010000  2.905000 4.165000 3.075000 ;
      RECT 3.155000  1.120000 3.530000 1.130000 ;
      RECT 3.155000  1.300000 3.530000 1.450000 ;
      RECT 3.155000  1.450000 3.325000 1.970000 ;
      RECT 3.325000  0.360000 4.225000 0.610000 ;
      RECT 3.350000  2.405000 3.665000 2.735000 ;
      RECT 3.495000  1.710000 5.060000 1.880000 ;
      RECT 3.495000  1.880000 3.665000 2.405000 ;
      RECT 3.715000  0.950000 3.885000 1.225000 ;
      RECT 3.715000  1.225000 4.130000 1.540000 ;
      RECT 3.835000  2.050000 4.165000 2.905000 ;
      RECT 4.055000  0.610000 4.225000 0.885000 ;
      RECT 4.055000  0.885000 4.470000 1.055000 ;
      RECT 4.300000  1.055000 4.470000 1.710000 ;
      RECT 4.375000  2.050000 5.640000 2.240000 ;
      RECT 4.375000  2.240000 6.955000 2.350000 ;
      RECT 4.395000  0.085000 4.645000 0.715000 ;
      RECT 4.525000  2.650000 5.140000 3.245000 ;
      RECT 4.735000  1.350000 5.060000 1.710000 ;
      RECT 4.875000  0.350000 5.400000 1.130000 ;
      RECT 5.230000  1.130000 5.400000 1.820000 ;
      RECT 5.230000  1.820000 5.640000 2.050000 ;
      RECT 5.310000  2.350000 6.955000 2.410000 ;
      RECT 5.310000  2.410000 5.640000 2.980000 ;
      RECT 5.695000  0.085000 6.025000 1.010000 ;
      RECT 5.810000  2.580000 6.140000 3.245000 ;
      RECT 6.625000  1.320000 6.955000 1.650000 ;
      RECT 6.710000  2.580000 7.040000 3.245000 ;
      RECT 6.785000  0.085000 7.045000 1.050000 ;
      RECT 6.785000  1.650000 6.955000 2.240000 ;
      RECT 7.215000  0.350000 7.545000 1.220000 ;
      RECT 7.215000  1.220000 8.230000 1.550000 ;
      RECT 7.215000  1.550000 7.545000 2.860000 ;
      RECT 7.775000  0.085000 8.035000 1.050000 ;
      RECT 7.775000  1.820000 8.025000 3.245000 ;
      RECT 8.745000  0.085000 9.005000 1.130000 ;
      RECT 8.755000  1.820000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_ls__dlrbn_2
END LIBRARY
