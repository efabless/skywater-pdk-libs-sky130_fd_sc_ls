# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__and3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.615000 1.450000 5.285000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.325000 4.335000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 3.230000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.350000 0.890000 0.960000 ;
        RECT 0.560000 0.960000 1.740000 1.130000 ;
        RECT 0.560000 1.130000 0.835000 1.800000 ;
        RECT 0.560000 1.800000 1.895000 1.970000 ;
        RECT 0.560000 1.970000 0.895000 2.980000 ;
        RECT 1.490000 0.350000 1.740000 0.960000 ;
        RECT 1.565000 1.970000 1.895000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 1.130000 ;
      RECT 1.035000  1.300000 2.235000 1.630000 ;
      RECT 1.065000  2.140000 1.395000 3.245000 ;
      RECT 1.070000  0.085000 1.320000 0.790000 ;
      RECT 1.920000  0.085000 2.250000 1.030000 ;
      RECT 2.065000  1.630000 2.235000 1.950000 ;
      RECT 2.065000  1.950000 5.625000 2.120000 ;
      RECT 2.065000  2.290000 2.395000 3.245000 ;
      RECT 2.420000  0.350000 2.670000 0.985000 ;
      RECT 2.420000  0.985000 4.090000 1.155000 ;
      RECT 2.565000  2.120000 2.895000 2.980000 ;
      RECT 2.850000  0.085000 3.180000 0.815000 ;
      RECT 3.065000  2.290000 3.645000 3.245000 ;
      RECT 3.410000  0.255000 5.640000 0.425000 ;
      RECT 3.410000  0.425000 3.740000 0.815000 ;
      RECT 3.815000  2.120000 4.145000 2.980000 ;
      RECT 3.920000  0.595000 4.090000 0.985000 ;
      RECT 4.310000  0.425000 4.640000 1.030000 ;
      RECT 4.315000  2.290000 4.645000 3.245000 ;
      RECT 4.810000  0.595000 5.140000 1.110000 ;
      RECT 4.810000  1.110000 5.625000 1.280000 ;
      RECT 4.815000  2.120000 5.145000 2.980000 ;
      RECT 5.310000  0.425000 5.640000 0.940000 ;
      RECT 5.315000  2.290000 5.645000 3.245000 ;
      RECT 5.455000  1.280000 5.625000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ls__and3_4
END LIBRARY
