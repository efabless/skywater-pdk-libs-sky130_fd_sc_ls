# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ls__a211o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.450000 6.115000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 0.255000 5.320000 0.505000 ;
        RECT 4.925000 0.505000 5.125000 0.670000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.470000 3.105000 1.720000 ;
        RECT 2.785000 1.720000 4.515000 1.890000 ;
        RECT 3.965000 1.470000 4.515000 1.720000 ;
        RECT 3.995000 1.890000 4.195000 2.150000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.450000 1.210000 3.780000 1.550000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.675000 1.240000 1.795000 1.410000 ;
        RECT 0.675000 1.410000 0.925000 1.720000 ;
        RECT 0.675000 1.720000 1.905000 1.890000 ;
        RECT 0.675000 1.890000 0.925000 2.980000 ;
        RECT 1.330000 0.350000 1.500000 0.790000 ;
        RECT 1.330000 0.790000 2.370000 0.960000 ;
        RECT 1.330000 0.960000 1.795000 1.240000 ;
        RECT 1.575000 1.890000 1.905000 2.980000 ;
        RECT 2.180000 0.545000 2.370000 0.790000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.225000  1.820000 0.475000 3.245000 ;
      RECT 0.820000  0.085000 1.150000 1.050000 ;
      RECT 1.125000  2.060000 1.375000 3.245000 ;
      RECT 1.680000  0.085000 2.010000 0.620000 ;
      RECT 1.965000  1.130000 3.280000 1.300000 ;
      RECT 1.965000  1.300000 2.615000 1.550000 ;
      RECT 2.105000  1.820000 2.275000 3.245000 ;
      RECT 2.445000  1.550000 2.615000 2.060000 ;
      RECT 2.445000  2.060000 3.825000 2.230000 ;
      RECT 2.540000  0.085000 2.870000 0.960000 ;
      RECT 2.545000  2.400000 4.710000 2.570000 ;
      RECT 2.545000  2.570000 2.875000 2.780000 ;
      RECT 3.040000  0.450000 3.280000 0.870000 ;
      RECT 3.040000  0.870000 4.245000 1.040000 ;
      RECT 3.040000  1.040000 3.280000 1.130000 ;
      RECT 3.045000  2.740000 4.300000 2.990000 ;
      RECT 3.460000  0.085000 3.790000 0.700000 ;
      RECT 3.960000  0.595000 4.245000 0.870000 ;
      RECT 3.960000  1.040000 4.245000 1.110000 ;
      RECT 3.960000  1.110000 6.055000 1.280000 ;
      RECT 4.420000  2.060000 6.910000 2.120000 ;
      RECT 4.420000  2.120000 5.960000 2.230000 ;
      RECT 4.420000  2.230000 4.710000 2.400000 ;
      RECT 4.425000  0.085000 4.755000 0.940000 ;
      RECT 4.500000  2.570000 4.710000 2.990000 ;
      RECT 4.880000  2.400000 5.555000 3.245000 ;
      RECT 5.295000  0.675000 6.405000 0.845000 ;
      RECT 5.680000  1.950000 6.910000 2.060000 ;
      RECT 5.725000  1.015000 6.055000 1.110000 ;
      RECT 5.725000  2.230000 5.960000 2.980000 ;
      RECT 6.130000  2.290000 6.460000 3.245000 ;
      RECT 6.235000  0.595000 6.405000 0.675000 ;
      RECT 6.235000  0.845000 6.405000 1.275000 ;
      RECT 6.580000  1.940000 6.910000 1.950000 ;
      RECT 6.585000  0.085000 6.915000 1.275000 ;
      RECT 6.630000  2.120000 6.910000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_ls__a211o_4
END LIBRARY
